module ALU #(
    parameter WIDTH = 32
) (
    ports
);
    
endmodule