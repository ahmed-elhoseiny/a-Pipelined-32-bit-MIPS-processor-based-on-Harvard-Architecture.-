module Hazard_Unit #(
parameter =,
) (

);
    
endmodule