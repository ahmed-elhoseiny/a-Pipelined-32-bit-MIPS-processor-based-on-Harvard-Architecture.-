module Fetch_stage #(
parameter
) (

);
    
endmodule